library ieee;
use ieee.std_logic_1164.all;

entity eightBitShifter_tb is
end eightBitShifter_tb;

architecture behav of eightBitShifter_tb is
component eightBitShifter
port(	i_e:	in std_logic_vector (7 downto 0);
	i_shift_in_e:	in std_logic;
	sel_e:	in std_logic_vector (1 downto 0);
	clock_e:	in std_logic;
	enable_e: in std_logic;
	clear_e: in std_logic;
	output_e:	out std_logic_vector (7 downto 0)
);
end component;


signal I, Output : std_logic_vector(7 downto 0);
signal I_SHIFT_IN, Clock, Enable, Clear : std_logic;
signal Sel : std_logic_vector(1 downto 0);

begin
eightBitShifter1: eightBitShifter port map (i_e => I, i_shift_in_e => I_SHIFT_IN, sel_e => Sel, clock_e => Clock, enable_e => Enable, clear_e => Clear, output_e => Output);

process
type pattern_type is record
I: std_logic_vector (7 downto 0);
I_SHIFT_IN, Clock, Enable, Clear: std_logic;
Sel: std_logic_vector(1 downto 0);
Output: std_logic_vector (7 downto 0);
end record;

type pattern_array is array (natural range <>) of pattern_type;
constant patterns : pattern_array :=
(("00000000", '0', '0', '1', '1', "11", "UUUUUUUU"), --initialization
("00000001", '1', '1', '1', '1', "11", "00000000"),
("00000001", '0', '0', '0', '0', "11", "00000000"),
("00000001", '1', '0', '0', '0', "11", "00000000"),
("00000001", '0', '1', '0', '0', "11", "00000000"),
("00000001", '0', '0', '1', '0', "11", "00000000"),
("00000001", '0', '0', '0', '1', "11", "00000000"),
("00000001", '1', '1', '0', '0', "11", "00000000"),
("00000001", '1', '0', '1', '0', "11", "00000000"),
("00000001", '1', '0', '0', '1', "11", "00000000"),
("00000001", '0', '1', '1', '0', "11", "00000001"),
("00000001", '0', '1', '0', '1', "11", "00000001"),
("00000001", '0', '0', '1', '1', "11", "00000001"),
("00000001", '1', '1', '1', '0', "11", "00000001"),
("00000001", '1', '1', '0', '1', "11", "00000001"),
("00000001", '1', '0', '1', '1', "11", "00000001"),
("00000001", '0', '1', '1', '1', "11", "00000000"),
("00000001", '1', '1', '1', '1', "10", "00000000"),
("00000001", '0', '0', '0', '0', "10", "00000000"),
("00000001", '1', '0', '0', '0', "10", "00000000"),
("00000001", '0', '1', '0', '0', "10", "00000000"),
("00000001", '0', '0', '1', '0', "10", "00000000"),
("00000001", '0', '0', '0', '1', "10", "00000000"),
("00000001", '1', '1', '0', '0', "10", "00000000"),
("00000001", '1', '0', '1', '0', "10", "00000000"),
("00000001", '1', '0', '0', '1', "10", "00000000"),
("00000001", '0', '1', '1', '0', "10", "00000000"),
("00000001", '0', '1', '0', '1', "10", "00000000"),
("00000001", '0', '0', '1', '1', "10", "00000000"),
("00000001", '1', '1', '1', '0', "10", "10000000"),
("00000001", '1', '1', '0', '1', "10", "10000000"),
("00000001", '1', '0', '1', '1', "10", "10000000"),
("00000001", '0', '1', '1', '1', "10", "00000000"),
("00000001", '1', '1', '1', '1', "01", "00000000"),
("00000001", '0', '0', '0', '0', "01", "00000000"),
("00000001", '1', '0', '0', '0', "01", "00000000"),
("00000001", '0', '1', '0', '0', "01", "00000000"),
("00000001", '0', '0', '1', '0', "01", "00000000"),
("00000001", '0', '0', '0', '1', "01", "00000000"),
("00000001", '1', '1', '0', '0', "01", "00000000"),
("00000001", '1', '0', '1', '0', "01", "00000000"),
("00000001", '1', '0', '0', '1', "01", "00000000"),
("00000001", '0', '1', '1', '0', "01", "00000010"),
("00000001", '0', '1', '0', '1', "01", "00000010"),
("00000001", '0', '0', '1', '1', "01", "00000010"),
("00000001", '1', '1', '1', '0', "01", "00000011"),
("00000001", '1', '1', '0', '1', "01", "00000011"),
("00000001", '1', '0', '1', '1', "01", "00000011"),
("00000001", '0', '1', '1', '1', "01", "00000000"),
("00000001", '1', '1', '1', '1', "00", "00000000"),
("00000001", '0', '0', '0', '0', "00", "00000000"),
("00000001", '1', '0', '0', '0', "00", "00000000"),
("00000001", '0', '1', '0', '0', "00", "00000000"),
("00000001", '0', '0', '1', '0', "00", "00000000"),
("00000001", '0', '0', '0', '1', "00", "00000000"),
("00000001", '1', '1', '0', '0', "00", "00000000"),
("00000001", '1', '0', '1', '0', "00", "00000000"),
("00000001", '1', '0', '0', '1', "00", "00000000"),
("00000001", '0', '1', '1', '0', "00", "00000000"),
("00000001", '0', '1', '0', '1', "00", "00000000"),
("00000001", '0', '0', '1', '1', "00", "00000000"),
("00000001", '1', '1', '1', '0', "00", "00000000"),
("00000001", '1', '1', '0', '1', "00", "00000000"),
("00000001", '1', '0', '1', '1', "00", "00000000"),
("00000001", '0', '1', '1', '1', "00", "00000000"));
begin

for n in patterns'range loop
I <= patterns(n).I;
I_SHIFT_IN <= patterns(n).I_SHIFT_IN;
Sel <= patterns(n).Sel;
Clock <= patterns(n).Clock;
Enable <= patterns(n).Enable;
Clear <= patterns(n).Clear;
wait for 1 ns;
assert Output = patterns(n).Output report (integer'image(n)) severity error;
if (n = 26 or n = 42) then
end if;
end loop;
assert false report "end of test" severity note;
wait;
end process;
end behav;
